module controller(
    input clk,
    input rst_n,
    input button,

    output save_A,
    output save_B,
    output show_result
);

    

endmodule