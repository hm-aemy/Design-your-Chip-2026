module controller(
    input logic clk,
    input logic rst_n,
    input logic button,

    output logic save_A,
    output logic save_B,
    output logic show_result
);



endmodule