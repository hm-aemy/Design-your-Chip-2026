module adder(
    input clk,
    input [3:0] operand,
    input save_A,
    input save_B,
    output [4:0] result
);

endmodule
