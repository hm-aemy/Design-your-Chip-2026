module seven_segment(
    input [3:0] digit,
    input update,
    output [6:0] seg
);

endmodule