module bcd_converter(
    input [4:0] binary,
    output [3:0] tens,
    output [3:0] ones
);

endmodule