module seven_segment(
    input logic        clk,
    input logic [3:0]  digit,
    input logic        update,
    output logic [6:0] seg
);

endmodule